`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Brandon Jamjampour
// Create date: 9/14/22 8:11pm
// description: behavior of norGATE
//////////////////////////////////////////////////////////////////////////////////


module NOR_GATE(
    input A,
    input B,
    output C
    );
    nor(C, B, A);
endmodule
