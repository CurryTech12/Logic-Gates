`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Engineer: Brandon Jamjampour
// Create Date: 09/14/2022 7:00pm
// Description: behavior of andGate

//////////////////////////////////////////////////////////////////////////////////


module AND_GATE(
    input A,
    input B,
    output C
    );
    and(C, B, A);
endmodule
