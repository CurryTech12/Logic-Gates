`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer:Brandon Jamjampour 
// desciprtion: behavior of a notGATE
// Create Date: 09/12/2022 8:00 PM
//////////////////////////////////////////////////////////////////////////////////


module NOT_GATE(
    input A,
    output B
    );
    not(B , A);
endmodule
