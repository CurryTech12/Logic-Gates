`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Brandon Jamjampour
// Create Date: 9/14/22 7:50pm
// Description: behavior of nandGATE

//////////////////////////////////////////////////////////////////////////////////


module NAND_GATE(
    input A,
    input B,
    output C
    );
    nand(C, B, A);
endmodule
