`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Engineer: Brandon Jamjampour
// Create Date: 9/14/22 7:32pm
// description: Time diagram of orGATE

//////////////////////////////////////////////////////////////////////////////////


module Or_GATE_(
    input A,
    input B,
    output C
    );
    or(C, B, A);
endmodule
