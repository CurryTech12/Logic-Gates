`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Engineer: Brandon Jamjampour
//Create date: 9/12/22 7:22pm
// description: behavior of xnorGATE
//////////////////////////////////////////////////////////////////////////////////


module XNOR_GATE(
    input A,
    input B,
    output C
    );
    xnor(C, B, A);
endmodule
